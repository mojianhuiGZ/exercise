module bus_arbiter;


endmodule
